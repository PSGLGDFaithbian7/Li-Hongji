`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/15 18:29:33
// Design Name: 
// Module Name: alu_eu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_eu(
input        rstn,
input [15:0] i_driveFromIssue_16,
output[15:0] o_freeToIssue_16,
//input [3:0]  i_controlFromIssue_4[15:0],//�����ź�
input [3:0]  i_controlFromIssue0_4,
input [3:0]  i_controlFromIssue1_4,
input [3:0]  i_controlFromIssue2_4,
input [3:0]  i_controlFromIssue3_4,
input [3:0]  i_controlFromIssue4_4,
input [3:0]  i_controlFromIssue5_4,
input [3:0]  i_controlFromIssue6_4,
input [3:0]  i_controlFromIssue7_4,
input [3:0]  i_controlFromIssue8_4,
input [3:0]  i_controlFromIssue9_4,
input [3:0]  i_controlFromIssue10_4,
input [3:0]  i_controlFromIssue11_4,
input [3:0]  i_controlFromIssue12_4,
input [3:0]  i_controlFromIssue13_4,
input [3:0]  i_controlFromIssue14_4,
input [3:0]  i_controlFromIssue15_4,
//input [3:0]  i_tagFromIssue_5[15:0],//ָ����
input [3:0]  i_tagFromIssue0_4,
input [3:0]  i_tagFromIssue1_4,
input [3:0]  i_tagFromIssue2_4,
input [3:0]  i_tagFromIssue3_4,
input [3:0]  i_tagFromIssue4_4,
input [3:0]  i_tagFromIssue5_4,
input [3:0]  i_tagFromIssue6_4,
input [3:0]  i_tagFromIssue7_4,
input [3:0]  i_tagFromIssue8_4,
input [3:0]  i_tagFromIssue9_4,
input [3:0]  i_tagFromIssue10_4,
input [3:0]  i_tagFromIssue11_4,
input [3:0]  i_tagFromIssue12_4,
input [3:0]  i_tagFromIssue13_4,
input [3:0]  i_tagFromIssue14_4,
input [3:0]  i_tagFromIssue15_4,
//input  [31:0] i_oprand1FromIssue_32[15:0],
input  [31:0] i_oprand1FromIssue0_32,
input  [31:0] i_oprand1FromIssue1_32,
input  [31:0] i_oprand1FromIssue2_32,
input  [31:0] i_oprand1FromIssue3_32,
input  [31:0] i_oprand1FromIssue4_32,
input  [31:0] i_oprand1FromIssue5_32,
input  [31:0] i_oprand1FromIssue6_32,
input  [31:0] i_oprand1FromIssue7_32,
input  [31:0] i_oprand1FromIssue8_32,
input  [31:0] i_oprand1FromIssue9_32,
input  [31:0] i_oprand1FromIssue10_32,
input  [31:0] i_oprand1FromIssue11_32,
input  [31:0] i_oprand1FromIssue12_32,
input  [31:0] i_oprand1FromIssue13_32,
input  [31:0] i_oprand1FromIssue14_32,
input  [31:0] i_oprand1FromIssue15_32,
//input  [31:0] i_oprand2FromIssue_32[15:0],
input  [31:0] i_oprand2FromIssue0_32,
input  [31:0] i_oprand2FromIssue1_32,
input  [31:0] i_oprand2FromIssue2_32,
input  [31:0] i_oprand2FromIssue3_32,
input  [31:0] i_oprand2FromIssue4_32,
input  [31:0] i_oprand2FromIssue5_32,
input  [31:0] i_oprand2FromIssue6_32,
input  [31:0] i_oprand2FromIssue7_32,
input  [31:0] i_oprand2FromIssue8_32,
input  [31:0] i_oprand2FromIssue9_32,
input  [31:0] i_oprand2FromIssue10_32,
input  [31:0] i_oprand2FromIssue11_32,
input  [31:0] i_oprand2FromIssue12_32,
input  [31:0] i_oprand2FromIssue13_32,
input  [31:0] i_oprand2FromIssue14_32,
input  [31:0] i_oprand2FromIssue15_32,
//input  [4:0]  i_areg_5[15:0],
input  [4:0]  i_areg0_5,
input  [4:0]  i_areg1_5,
input  [4:0]  i_areg2_5,
input  [4:0]  i_areg3_5,
input  [4:0]  i_areg4_5,
input  [4:0]  i_areg5_5,
input  [4:0]  i_areg6_5,
input  [4:0]  i_areg7_5,
input  [4:0]  i_areg8_5,
input  [4:0]  i_areg9_5,
input  [4:0]  i_areg10_5,
input  [4:0]  i_areg11_5,
input  [4:0]  i_areg12_5,
input  [4:0]  i_areg13_5,
input  [4:0]  i_areg14_5,
input  [4:0]  i_areg15_5,

output[15:0] o_driveToIssue_16,
input [15:0] i_freeFromIssue_16,
//output [31:0] o_resultToIssue_32[15:0],
output [31:0] o_resultToIssue0_32,
output [31:0] o_resultToIssue1_32,
output [31:0] o_resultToIssue2_32,
output [31:0] o_resultToIssue3_32,
output [31:0] o_resultToIssue4_32,
output [31:0] o_resultToIssue5_32,
output [31:0] o_resultToIssue6_32,
output [31:0] o_resultToIssue7_32,
output [31:0] o_resultToIssue8_32,
output [31:0] o_resultToIssue9_32,
output [31:0] o_resultToIssue10_32,
output [31:0] o_resultToIssue11_32,
output [31:0] o_resultToIssue12_32,
output [31:0] o_resultToIssue13_32,
output [31:0] o_resultToIssue14_32,
output [31:0] o_resultToIssue15_32,
//output [3:0]  o_indexToIssue_4[15:0],
output [3:0]  o_indexToIssue0_4,
output [3:0]  o_indexToIssue1_4,
output [3:0]  o_indexToIssue2_4,
output [3:0]  o_indexToIssue3_4,
output [3:0]  o_indexToIssue4_4,
output [3:0]  o_indexToIssue5_4,
output [3:0]  o_indexToIssue6_4,
output [3:0]  o_indexToIssue7_4,
output [3:0]  o_indexToIssue8_4,
output [3:0]  o_indexToIssue9_4,
output [3:0]  o_indexToIssue10_4,
output [3:0]  o_indexToIssue11_4,
output [3:0]  o_indexToIssue12_4,
output [3:0]  o_indexToIssue13_4,
output [3:0]  o_indexToIssue14_4,
output [3:0]  o_indexToIssue15_4,
output[15:0] o_driveToMD_16,
input [15:0] i_freeFromMD_16,
//output [31:0]o_resultToMD_32[15:0],
output [31:0]o_resultToMD0_32,
output [31:0]o_resultToMD1_32,
output [31:0]o_resultToMD2_32,
output [31:0]o_resultToMD3_32,
output [31:0]o_resultToMD4_32,
output [31:0]o_resultToMD5_32,
output [31:0]o_resultToMD6_32,
output [31:0]o_resultToMD7_32,
output [31:0]o_resultToMD8_32,
output [31:0]o_resultToMD9_32,
output [31:0]o_resultToMD10_32,
output [31:0]o_resultToMD11_32,
output [31:0]o_resultToMD12_32,
output [31:0]o_resultToMD13_32,
output [31:0]o_resultToMD14_32,
output [31:0]o_resultToMD15_32,
//output [3:0] o_indexToMD_4[15:0],
output [3:0] o_indexToMD0_4,
output [3:0] o_indexToMD1_4,
output [3:0] o_indexToMD2_4,
output [3:0] o_indexToMD3_4,
output [3:0] o_indexToMD4_4,
output [3:0] o_indexToMD5_4,
output [3:0] o_indexToMD6_4,
output [3:0] o_indexToMD7_4,
output [3:0] o_indexToMD8_4,
output [3:0] o_indexToMD9_4,
output [3:0] o_indexToMD10_4,
output [3:0] o_indexToMD11_4,
output [3:0] o_indexToMD12_4,
output [3:0] o_indexToMD13_4,
output [3:0] o_indexToMD14_4,
output [3:0] o_indexToMD15_4,
output[15:0] o_driveToBranch_16,
input [15:0] i_freeFromBranch_16,
//output  [31:0]o_resultToBranch_32[15:0],
output  [31:0]o_resultToBranch0_32,
output  [31:0]o_resultToBranch1_32,
output  [31:0]o_resultToBranch2_32,
output  [31:0]o_resultToBranch3_32,
output  [31:0]o_resultToBranch4_32,
output  [31:0]o_resultToBranch5_32,
output  [31:0]o_resultToBranch6_32,
output  [31:0]o_resultToBranch7_32,
output  [31:0]o_resultToBranch8_32,
output  [31:0]o_resultToBranch9_32,
output  [31:0]o_resultToBranch10_32,
output  [31:0]o_resultToBranch11_32,
output  [31:0]o_resultToBranch12_32,
output  [31:0]o_resultToBranch13_32,
output  [31:0]o_resultToBranch14_32,
output  [31:0]o_resultToBranch15_32,
//output  [3:0] o_indexToBranch_4[15:0],
output  [3:0] o_indexToBranch0_4,
output  [3:0] o_indexToBranch1_4,
output  [3:0] o_indexToBranch2_4,
output  [3:0] o_indexToBranch3_4,
output  [3:0] o_indexToBranch4_4,
output  [3:0] o_indexToBranch5_4,
output  [3:0] o_indexToBranch6_4,
output  [3:0] o_indexToBranch7_4,
output  [3:0] o_indexToBranch8_4,
output  [3:0] o_indexToBranch9_4,
output  [3:0] o_indexToBranch10_4,
output  [3:0] o_indexToBranch11_4,
output  [3:0] o_indexToBranch12_4,
output  [3:0] o_indexToBranch13_4,
output  [3:0] o_indexToBranch14_4,
output  [3:0] o_indexToBranch15_4,
output[15:0] o_driveToWB_16,
input [15:0] i_freeFromWB_16,
//output [31:0]o_resultToWB_32[15:0],
output [31:0]o_resultToWB0_32,
output [31:0]o_resultToWB1_32,
output [31:0]o_resultToWB2_32,
output [31:0]o_resultToWB3_32,
output [31:0]o_resultToWB4_32,
output [31:0]o_resultToWB5_32,
output [31:0]o_resultToWB6_32,
output [31:0]o_resultToWB7_32,
output [31:0]o_resultToWB8_32,
output [31:0]o_resultToWB9_32,
output [31:0]o_resultToWB10_32,
output [31:0]o_resultToWB11_32,
output [31:0]o_resultToWB12_32,
output [31:0]o_resultToWB13_32,
output [31:0]o_resultToWB14_32,
output [31:0]o_resultToWB15_32,
output [15:0]o_indexToWB_16,
//output [4:0]  o_areg_5[15:0]
output [4:0]  o_areg0_5,
output [4:0]  o_areg1_5,
output [4:0]  o_areg2_5,
output [4:0]  o_areg3_5,
output [4:0]  o_areg4_5,
output [4:0]  o_areg5_5,
output [4:0]  o_areg6_5,
output [4:0]  o_areg7_5,
output [4:0]  o_areg8_5,
output [4:0]  o_areg9_5,
output [4:0]  o_areg10_5,
output [4:0]  o_areg11_5,
output [4:0]  o_areg12_5,
output [4:0]  o_areg13_5,
output [4:0]  o_areg14_5,
output [4:0]  o_areg15_5
    );
     alu  alu0(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[0]),
             .o_freeToIssue(o_freeToIssue_16[0]),
             .i_controlFromIssue_4(i_controlFromIssue0_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue0_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue0_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue0_32),
             .i_areg_5(i_areg0_5),

             .o_driveToIssue(o_driveToIssue_16[0]),
             .i_freeFromIssue(i_freeFromIssue_16[0]),
             .o_resultToIssue_32(o_resultToIssue0_32),
             .o_indexToIssue_4(o_indexToIssue0_4),
             .o_driveToMD(o_driveToMD_16[0]),
             .i_freeFromMD(i_freeFromMD_16[0]),
             .o_resultToMD_32(o_resultToMD0_32),
             .o_indexToMD_4(o_indexToMD0_4),
             .o_driveToBranch(o_driveToBranch_16[0]),
             .i_freeFromBranch(i_freeFromBranch_16[0]),
             .o_resultToBranch_32(o_resultToBranch0_32),
             .o_indexToBranch_4(o_indexToBranch0_4),
             .o_driveToWB(o_driveToWB_16[0]),
             .i_freeFromWB(i_freeFromWB_16[0]),
             .o_resultToWB_32(o_resultToWB0_32),
             .o_indexToWB(o_indexToWB_16[0]),
             .o_areg_5(o_areg0_5)
                );
    alu  alu1(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[1]),
             .o_freeToIssue(o_freeToIssue_16[1]),
             .i_controlFromIssue_4(i_controlFromIssue1_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue1_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue1_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue1_32),
             .i_areg_5(i_areg1_5),

             .o_driveToIssue(o_driveToIssue_16[1]),
             .i_freeFromIssue(i_freeFromIssue_16[1]),
             .o_resultToIssue_32(o_resultToIssue1_32),
             .o_indexToIssue_4(o_indexToIssue1_4),
             .o_driveToMD(o_driveToMD_16[1]),
             .i_freeFromMD(i_freeFromMD_16[1]),
             .o_resultToMD_32(o_resultToMD1_32),
             .o_indexToMD_4(o_indexToMD1_4),
             .o_driveToBranch(o_driveToBranch_16[1]),
             .i_freeFromBranch(i_freeFromBranch_16[1]),
             .o_resultToBranch_32(o_resultToBranch1_32),
             .o_indexToBranch_4(o_indexToBranch1_4),
             .o_driveToWB(o_driveToWB_16[1]),
             .i_freeFromWB(i_freeFromWB_16[1]),
             .o_resultToWB_32(o_resultToWB1_32),
             .o_indexToWB(o_indexToWB_16[1]),
             .o_areg_5(o_areg1_5)
      );
      alu  alu2(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[2]),
             .o_freeToIssue(o_freeToIssue_16[2]),
             .i_controlFromIssue_4(i_controlFromIssue2_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue2_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue2_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue2_32),
             .i_areg_5(i_areg2_5),

             .o_driveToIssue(o_driveToIssue_16[2]),
             .i_freeFromIssue(i_freeFromIssue_16[2]),
             .o_resultToIssue_32(o_resultToIssue2_32),
             .o_indexToIssue_4(o_indexToIssue2_4),
             .o_driveToMD(o_driveToMD_16[2]),
             .i_freeFromMD(i_freeFromMD_16[2]),
             .o_resultToMD_32(o_resultToMD2_32),
             .o_indexToMD_4(o_indexToMD2_4),
             .o_driveToBranch(o_driveToBranch_16[2]),
             .i_freeFromBranch(i_freeFromBranch_16[2]),
             .o_resultToBranch_32(o_resultToBranch2_32),
             .o_indexToBranch_4(o_indexToBranch2_4),
             .o_driveToWB(o_driveToWB_16[2]),
             .i_freeFromWB(i_freeFromWB_16[2]),
             .o_resultToWB_32(o_resultToWB2_32),
             .o_indexToWB(o_indexToWB_16[2]),
             .o_areg_5(o_areg2_5)
     );
      alu  alu3(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[3]),
             .o_freeToIssue(o_freeToIssue_16[3]),
             .i_controlFromIssue_4(i_controlFromIssue3_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue3_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue3_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue3_32),
             .i_areg_5(i_areg3_5),

             .o_driveToIssue(o_driveToIssue_16[3]),
             .i_freeFromIssue(i_freeFromIssue_16[3]),
             .o_resultToIssue_32(o_resultToIssue3_32),
             .o_indexToIssue_4(o_indexToIssue3_4),
             .o_driveToMD(o_driveToMD_16[3]),
             .i_freeFromMD(i_freeFromMD_16[3]),
             .o_resultToMD_32(o_resultToMD3_32),
             .o_indexToMD_4(o_indexToMD3_4),
             .o_driveToBranch(o_driveToBranch_16[3]),
             .i_freeFromBranch(i_freeFromBranch_16[3]),
             .o_resultToBranch_32(o_resultToBranch3_32),
             .o_indexToBranch_4(o_indexToBranch3_4),
             .o_driveToWB(o_driveToWB_16[3]),
             .i_freeFromWB(i_freeFromWB_16[3]),
             .o_resultToWB_32(o_resultToWB3_32),
             .o_indexToWB(o_indexToWB_16[3]),
             .o_areg_5(o_areg3_5)
     );
      alu  alu4(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[4]),
             .o_freeToIssue(o_freeToIssue_16[4]),
             .i_controlFromIssue_4(i_controlFromIssue4_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue4_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue4_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue4_32),
             .i_areg_5(i_areg4_5),

             .o_driveToIssue(o_driveToIssue_16[4]),
             .i_freeFromIssue(i_freeFromIssue_16[4]),
             .o_resultToIssue_32(o_resultToIssue4_32),
             .o_indexToIssue_4(o_indexToIssue4_4),
             .o_driveToMD(o_driveToMD_16[4]),
             .i_freeFromMD(i_freeFromMD_16[4]),
             .o_resultToMD_32(o_resultToMD4_32),
             .o_indexToMD_4(o_indexToMD4_4),
             .o_driveToBranch(o_driveToBranch_16[4]),
             .i_freeFromBranch(i_freeFromBranch_16[4]),
             .o_resultToBranch_32(o_resultToBranch4_32),
             .o_indexToBranch_4(o_indexToBranch4_4),
             .o_driveToWB(o_driveToWB_16[4]),
             .i_freeFromWB(i_freeFromWB_16[4]),
             .o_resultToWB_32(o_resultToWB4_32),
             .o_indexToWB(o_indexToWB_16[4]),
             .o_areg_5(o_areg4_5)
     );
      alu  alu5(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[5]),
             .o_freeToIssue(o_freeToIssue_16[5]),
             .i_controlFromIssue_4(i_controlFromIssue5_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue5_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue5_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue5_32),
             .i_areg_5(i_areg5_5),

             .o_driveToIssue(o_driveToIssue_16[5]),
             .i_freeFromIssue(i_freeFromIssue_16[5]),
             .o_resultToIssue_32(o_resultToIssue5_32),
             .o_indexToIssue_4(o_indexToIssue5_4),
             .o_driveToMD(o_driveToMD_16[5]),
             .i_freeFromMD(i_freeFromMD_16[5]),
             .o_resultToMD_32(o_resultToMD5_32),
             .o_indexToMD_4(o_indexToMD5_4),
             .o_driveToBranch(o_driveToBranch_16[5]),
             .i_freeFromBranch(i_freeFromBranch_16[5]),
             .o_resultToBranch_32(o_resultToBranch5_32),
             .o_indexToBranch_4(o_indexToBranch5_4),
             .o_driveToWB(o_driveToWB_16[5]),
             .i_freeFromWB(i_freeFromWB_16[5]),
             .o_resultToWB_32(o_resultToWB5_32),
             .o_indexToWB(o_indexToWB_16[5]),
             .o_areg_5(o_areg5_5)
     );
      alu  alu6(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[6]),
             .o_freeToIssue(o_freeToIssue_16[6]),
             .i_controlFromIssue_4(i_controlFromIssue6_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue6_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue6_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue6_32),
             .i_areg_5(i_areg6_5),

             .o_driveToIssue(o_driveToIssue_16[6]),
             .i_freeFromIssue(i_freeFromIssue_16[6]),
             .o_resultToIssue_32(o_resultToIssue6_32),
             .o_indexToIssue_4(o_indexToIssue6_4),
             .o_driveToMD(o_driveToMD_16[6]),
             .i_freeFromMD(i_freeFromMD_16[6]),
             .o_resultToMD_32(o_resultToMD6_32),
             .o_indexToMD_4(o_indexToMD6_4),
             .o_driveToBranch(o_driveToBranch_16[6]),
             .i_freeFromBranch(i_freeFromBranch_16[6]),
             .o_resultToBranch_32(o_resultToBranch6_32),
             .o_indexToBranch_4(o_indexToBranch6_4),
             .o_driveToWB(o_driveToWB_16[6]),
             .i_freeFromWB(i_freeFromWB_16[6]),
             .o_resultToWB_32(o_resultToWB6_32),
             .o_indexToWB(o_indexToWB_16[6]),
             .o_areg_5(o_areg6_5)
     );
      alu  alu7(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[7]),
             .o_freeToIssue(o_freeToIssue_16[7]),
             .i_controlFromIssue_4(i_controlFromIssue7_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue7_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue7_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue7_32),
             .i_areg_5(i_areg7_5),

             .o_driveToIssue(o_driveToIssue_16[7]),
             .i_freeFromIssue(i_freeFromIssue_16[7]),
             .o_resultToIssue_32(o_resultToIssue7_32),
             .o_indexToIssue_4(o_indexToIssue7_4),
             .o_driveToMD(o_driveToMD_16[7]),
             .i_freeFromMD(i_freeFromMD_16[7]),
             .o_resultToMD_32(o_resultToMD7_32),
             .o_indexToMD_4(o_indexToMD7_4),
             .o_driveToBranch(o_driveToBranch_16[7]),
             .i_freeFromBranch(i_freeFromBranch_16[7]),
             .o_resultToBranch_32(o_resultToBranch7_32),
             .o_indexToBranch_4(o_indexToBranch7_4),
             .o_driveToWB(o_driveToWB_16[7]),
             .i_freeFromWB(i_freeFromWB_16[7]),
             .o_resultToWB_32(o_resultToWB7_32),
             .o_indexToWB(o_indexToWB_16[7]),
             .o_areg_5(o_areg7_5)
     );
      alu  alu8(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[8]),
             .o_freeToIssue(o_freeToIssue_16[8]),
             .i_controlFromIssue_4(i_controlFromIssue8_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue8_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue8_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue8_32),
             .i_areg_5(i_areg8_5),

             .o_driveToIssue(o_driveToIssue_16[8]),
             .i_freeFromIssue(i_freeFromIssue_16[8]),
             .o_resultToIssue_32(o_resultToIssue8_32),
             .o_indexToIssue_4(o_indexToIssue8_4),
             .o_driveToMD(o_driveToMD_16[8]),
             .i_freeFromMD(i_freeFromMD_16[8]),
             .o_resultToMD_32(o_resultToMD8_32),
             .o_indexToMD_4(o_indexToMD8_4),
             .o_driveToBranch(o_driveToBranch_16[8]),
             .i_freeFromBranch(i_freeFromBranch_16[8]),
             .o_resultToBranch_32(o_resultToBranch8_32),
             .o_indexToBranch_4(o_indexToBranch8_4),
             .o_driveToWB(o_driveToWB_16[8]),
             .i_freeFromWB(i_freeFromWB_16[8]),
             .o_resultToWB_32(o_resultToWB8_32),
             .o_indexToWB(o_indexToWB_16[8]),
             .o_areg_5(o_areg8_5)
     );
      alu  alu9(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[9]),
             .o_freeToIssue(o_freeToIssue_16[9]),
             .i_controlFromIssue_4(i_controlFromIssue9_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue9_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue9_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue9_32),
             .i_areg_5(i_areg9_5),

             .o_driveToIssue(o_driveToIssue_16[9]),
             .i_freeFromIssue(i_freeFromIssue_16[9]),
             .o_resultToIssue_32(o_resultToIssue9_32),
             .o_indexToIssue_4(o_indexToIssue9_4),
             .o_driveToMD(o_driveToMD_16[9]),
             .i_freeFromMD(i_freeFromMD_16[9]),
             .o_resultToMD_32(o_resultToMD9_32),
             .o_indexToMD_4(o_indexToMD9_4),
             .o_driveToBranch(o_driveToBranch_16[9]),
             .i_freeFromBranch(i_freeFromBranch_16[9]),
             .o_resultToBranch_32(o_resultToBranch9_32),
             .o_indexToBranch_4(o_indexToBranch9_4),
             .o_driveToWB(o_driveToWB_16[9]),
             .i_freeFromWB(i_freeFromWB_16[9]),
             .o_resultToWB_32(o_resultToWB9_32),
             .o_indexToWB(o_indexToWB_16[9]),
             .o_areg_5(o_areg9_5)
     );
      alu  alu10(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[10]),
             .o_freeToIssue(o_freeToIssue_16[10]),
             .i_controlFromIssue_4(i_controlFromIssue10_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue10_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue10_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue10_32),
             .i_areg_5(i_areg10_5),

             .o_driveToIssue(o_driveToIssue_16[10]),
             .i_freeFromIssue(i_freeFromIssue_16[10]),
             .o_resultToIssue_32(o_resultToIssue10_32),
             .o_indexToIssue_4(o_indexToIssue10_4),
             .o_driveToMD(o_driveToMD_16[10]),
             .i_freeFromMD(i_freeFromMD_16[10]),
             .o_resultToMD_32(o_resultToMD10_32),
             .o_indexToMD_4(o_indexToMD10_4),
             .o_driveToBranch(o_driveToBranch_16[10]),
             .i_freeFromBranch(i_freeFromBranch_16[10]),
             .o_resultToBranch_32(o_resultToBranch10_32),
             .o_indexToBranch_4(o_indexToBranch10_4),
             .o_driveToWB(o_driveToWB_16[10]),
             .i_freeFromWB(i_freeFromWB_16[10]),
             .o_resultToWB_32(o_resultToWB10_32),
             .o_indexToWB(o_indexToWB_16[10]),
             .o_areg_5(o_areg10_5)
     );
      alu  alu11(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[11]),
             .o_freeToIssue(o_freeToIssue_16[11]),
             .i_controlFromIssue_4(i_controlFromIssue11_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue11_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue11_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue11_32),
             .i_areg_5(i_areg11_5),

             .o_driveToIssue(o_driveToIssue_16[11]),
             .i_freeFromIssue(i_freeFromIssue_16[11]),
             .o_resultToIssue_32(o_resultToIssue11_32),
             .o_indexToIssue_4(o_indexToIssue11_4),
             .o_driveToMD(o_driveToMD_16[11]),
             .i_freeFromMD(i_freeFromMD_16[11]),
             .o_resultToMD_32(o_resultToMD11_32),
             .o_indexToMD_4(o_indexToMD11_4),
             .o_driveToBranch(o_driveToBranch_16[11]),
             .i_freeFromBranch(i_freeFromBranch_16[11]),
             .o_resultToBranch_32(o_resultToBranch11_32),
             .o_indexToBranch_4(o_indexToBranch11_4),
             .o_driveToWB(o_driveToWB_16[11]),
             .i_freeFromWB(i_freeFromWB_16[11]),
             .o_resultToWB_32(o_resultToWB11_32),
             .o_indexToWB(o_indexToWB_16[11]),
             .o_areg_5(o_areg11_5)
     );
      alu  alu12(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[12]),
             .o_freeToIssue(o_freeToIssue_16[12]),
             .i_controlFromIssue_4(i_controlFromIssue12_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue12_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue12_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue12_32),
             .i_areg_5(i_areg12_5),

             .o_driveToIssue(o_driveToIssue_16[12]),
             .i_freeFromIssue(i_freeFromIssue_16[12]),
             .o_resultToIssue_32(o_resultToIssue12_32),
             .o_indexToIssue_4(o_indexToIssue12_4),
             .o_driveToMD(o_driveToMD_16[12]),
             .i_freeFromMD(i_freeFromMD_16[12]),
             .o_resultToMD_32(o_resultToMD12_32),
             .o_indexToMD_4(o_indexToMD12_4),
             .o_driveToBranch(o_driveToBranch_16[12]),
             .i_freeFromBranch(i_freeFromBranch_16[12]),
             .o_resultToBranch_32(o_resultToBranch12_32),
             .o_indexToBranch_4(o_indexToBranch12_4),
             .o_driveToWB(o_driveToWB_16[12]),
             .i_freeFromWB(i_freeFromWB_16[12]),
             .o_resultToWB_32(o_resultToWB12_32),
             .o_indexToWB(o_indexToWB_16[12]),
             .o_areg_5(o_areg12_5)
     );
      alu  alu13(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[13]),
             .o_freeToIssue(o_freeToIssue_16[13]),
             .i_controlFromIssue_4(i_controlFromIssue13_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue13_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue13_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue13_32),
             .i_areg_5(i_areg13_5),

             .o_driveToIssue(o_driveToIssue_16[13]),
             .i_freeFromIssue(i_freeFromIssue_16[13]),
             .o_resultToIssue_32(o_resultToIssue13_32),
             .o_indexToIssue_4(o_indexToIssue13_4),
             .o_driveToMD(o_driveToMD_16[13]),
             .i_freeFromMD(i_freeFromMD_16[13]),
             .o_resultToMD_32(o_resultToMD13_32),
             .o_indexToMD_4(o_indexToMD13_4),
             .o_driveToBranch(o_driveToBranch_16[13]),
             .i_freeFromBranch(i_freeFromBranch_16[13]),
             .o_resultToBranch_32(o_resultToBranch13_32),
             .o_indexToBranch_4(o_indexToBranch13_4),
             .o_driveToWB(o_driveToWB_16[13]),
             .i_freeFromWB(i_freeFromWB_16[13]),
             .o_resultToWB_32(o_resultToWB13_32),
             .o_indexToWB(o_indexToWB_16[13]),
             .o_areg_5(o_areg13_5)
     );
     alu  alu14(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[14]),
             .o_freeToIssue(o_freeToIssue_16[14]),
             .i_controlFromIssue_4(i_controlFromIssue14_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue14_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue14_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue14_32),
             .i_areg_5(i_areg14_5),

             .o_driveToIssue(o_driveToIssue_16[14]),
             .i_freeFromIssue(i_freeFromIssue_16[14]),
             .o_resultToIssue_32(o_resultToIssue14_32),
             .o_indexToIssue_4(o_indexToIssue14_4),
             .o_driveToMD(o_driveToMD_16[14]),
             .i_freeFromMD(i_freeFromMD_16[14]),
             .o_resultToMD_32(o_resultToMD14_32),
             .o_indexToMD_4(o_indexToMD14_4),
             .o_driveToBranch(o_driveToBranch_16[14]),
             .i_freeFromBranch(i_freeFromBranch_16[14]),
             .o_resultToBranch_32(o_resultToBranch14_32),
             .o_indexToBranch_4(o_indexToBranch14_4),
             .o_driveToWB(o_driveToWB_16[14]),
             .i_freeFromWB(i_freeFromWB_16[14]),
             .o_resultToWB_32(o_resultToWB14_32),
             .o_indexToWB(o_indexToWB_16[14]),
             .o_areg_5(o_areg14_5)
     );
     alu  alu15(
             .rstn(rstn),
             .i_driveFromIssue(i_driveFromIssue_16[15]),
             .o_freeToIssue(o_freeToIssue_16[15]),
             .i_controlFromIssue_4(i_controlFromIssue15_4),//�����ź�
             .i_tagFromIssue_4(i_tagFromIssue15_4),//ָ����+��·��־λ
             .i_oprand1FromIssue_32(i_oprand1FromIssue15_32),
             .i_oprand2FromIssue_32(i_oprand2FromIssue15_32),
             .i_areg_5(i_areg15_5),

             .o_driveToIssue(o_driveToIssue_16[15]),
             .i_freeFromIssue(i_freeFromIssue_16[15]),
             .o_resultToIssue_32(o_resultToIssue15_32),
             .o_indexToIssue_4(o_indexToIssue15_4),
             .o_driveToMD(o_driveToMD_16[15]),
             .i_freeFromMD(i_freeFromMD_16[15]),
             .o_resultToMD_32(o_resultToMD15_32),
             .o_indexToMD_4(o_indexToMD15_4),
             .o_driveToBranch(o_driveToBranch_16[15]),
             .i_freeFromBranch(i_freeFromBranch_16[15]),
             .o_resultToBranch_32(o_resultToBranch15_32),
             .o_indexToBranch_4(o_indexToBranch15_4),
             .o_driveToWB(o_driveToWB_16[15]),
             .i_freeFromWB(i_freeFromWB_16[15]),
             .o_resultToWB_32(o_resultToWB15_32),
             .o_indexToWB(o_indexToWB_16[15]),
             .o_areg_5(o_areg15_5)
     );           
endmodule
